

class mem_model_base_test extends uvm_test;

  `uvm_component_utils(mem_model_base_test)

  // Environment class instantiation.
  mem_env env;

  // Environment configuration object instantiation.
  mem_env_config env_config;

  //---------------------------------------
  // constructor
  //---------------------------------------
  function new(string name = "mem_model_base_test",uvm_component parent=null);
    super.new(name,parent);
  endfunction : new

  //---------------------------------------
  // build_phase
  //---------------------------------------
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    // Create environment and its configuration object.
    env = mem_env::type_id::create("env", this);
    env_config = mem_env_config::type_id::create("env_config", this);

    // Configure Agent.
    env_config.mem_agent_cnfg = mem_agent_config::type_id::create("mem_agent_cnfg");
    env_config.mem_agent_cnfg.active = UVM_ACTIVE;

    // Post configure and set configuration object to database
    uvm_config_db#(mem_env_config)::set(uvm_root::get(), "*", "mem_env_config", env_config);

  endfunction : build_phase

  //---------------------------------------
  // end_of_elobaration phase
  //---------------------------------------
  virtual function void end_of_elaboration();
    //print's the topology
    print();
  endfunction

  //---------------------------------------
  // end_of_elobaration phase
  //---------------------------------------
 function void report_phase(uvm_phase phase);
   uvm_report_server svr;
   super.report_phase(phase);

   svr = uvm_report_server::get_server();
   if(svr.get_severity_count(UVM_FATAL)+svr.get_severity_count(UVM_ERROR)>0) begin
     `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
     `uvm_info(get_type_name(), "----            TEST FAIL          ----", UVM_NONE)
     `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
    end
    else begin
     `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
     `uvm_info(get_type_name(), "----           TEST PASS           ----", UVM_NONE)
     `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
    end
  endfunction

endclass : mem_model_base_test
