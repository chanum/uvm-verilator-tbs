
package mem_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "mem_seq_item.svh"
  // `include "mem_agent_config.svh"
  `include "mem_driver.svh"
  `include "mem_monitor.svh"
  `include "mem_sequencer.svh"
  `include "mem_agent.svh"

  // Utility sequences
  `include "mem_sequence.svh"

endpackage : mem_agent_pkg