
package ct_param_in_agent_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ct_param_in_seq_item.svh"
  `include "ct_param_in_agent_config.svh"
  `include "ct_param_in_driver.svh"
  `include "ct_param_in_monitor.svh"
  `include "ct_param_in_sequencer.svh"
  `include "ct_param_in_agent.svh"

  // Utility sequences
  // `include "ct_param_in_seq.svh"

endpackage